Hund

Från Wikipedia
För andra betydelser, se Hund (olika betydelser).
Hund

Norsk älghund, grå (gråhund)
Systematik
Domän	Eukaryoter
Eukaryota
Rike	Djur
Animalia
Stam	Ryggsträngsdjur
Chordata
Understam	Ryggradsdjur
Vertebrata
Klass	Däggdjur
Mammalia
Ordning	Rovdjur
Carnivora
Familj	Hunddjur
Canidae
Släkte	Canis
Art	Varg
Canis lupus
Underart	Hund
C. l. familiaris
Vetenskapligt namn
§Canis lupus familiaris
Auktor	Linné, 1758
Hitta fler artiklar om djur med
Djurportalen
Hund (Canis lupus familiaris eller Canis lupus domesticus, tidigare även Canis familiaris) är en domesticerad underart av varg (Canis lupus). Hundar finns av många olika raser, vilka i Sverige organiseras av Svenska Kennelklubben (SKK), riksorganisation för svenska hundägare. Den vetenskapliga läran om hundar kallas kynologi. En hund av hankön kallas hund[1] och en av honkön kallas för tik och dess avkomma kallas valp. Det finns cirka 800 000 hundar i Sverige varav drygt 500 000 är registrerade hos Svenska Kennelklubben.[2] Dessa är fördelade på cirka 600 000 hushåll[3].

Innehåll

1 Taxonomi
1.1 Släktskap mellan hundraser
2 Historia
3 Födoämnen, skötsel och vård
4 Fortplantning och avel
5 Hundens användningsområden
5.1 Familjehundar
5.2 Jakthundar
5.3 Brukshundar
5.4 Hundsport
5.5 Utställning
5.6 Draghund
6 Hundraser
6.1 Att välja en ras som passar
6.2 Valets kval
6.3 Allergivänliga raser
6.4 Svenska hundraser
6.5 Förbjudna hundraser
7 Övrigt och kuriosa
8 Galleri
9 Se även
10 Källor
11 Noter
12 Externa länkar
Taxonomi

Huruvida hunden är en underart, Canis lupus familiaris, till vargen (Canis lupus) har diskuterats eftersom detta medför att de hundraser som vi känner idag klassificeras som varianter och subvarianter. Detta gör att vissa forskare fortfarande vill hävda hunden som egen art, Canis familiaris, precis som Linné gjorde 1758, när han beskrev den. Senare forskning kring hundens DNA har dock påvisat hundens släktskap med vargen, och därför reklassificerade man den som en underart av varg 1993.

Släktskap mellan hundraser

En studie ledd av Elaine Ostrander, genetiker vid Fred Hutchinson Cancer Research Center vid University of Washington, har förändrat synen på ålder och släktskap bland hundraser.[4] Deras analyser av mitokondrie-DNA har bland annat visat att schäfer är närmare släkt med mastiff, boxer och andra typiska vakthundar än de fårhundar de vanligtvis klassificeras tillsammans med. Samma analyser visar också att raser som greyhound, irländsk varghund, borzoi och sanktbernhardshund bär släktskap med fårhund. Studien har vidare resulterat i att vissa rasers ålder har måst omvärderas. Raser som tidigare ansetts tillhöra de absolut äldsta som gråhund, faraohund och ibizahund kanske inte är äldre än 150–200 år gamla i nuvarande form.

Historia

Hunden är en av människans äldsta följeslagare. Hunden härstammar från domesticerade vargar, som antingen uppkommit genom att vargungar uppfostrats av människor, eller att vargflockar uppehållit sig kring mänskliga boplatser, där de levde på människans matrester och blivit tamare för varje generation. Det finns kvarlevor från hund i människans sällskap i Östasien möjligen från 30 000 fvt och med största säkerhet 7 000 fvt, bl.a. de s.k. torvhundarna. Nya forskningsrön (2011) från KTH bekräftar att Asien söder om Yangtzefloden var den viktigaste och kanske enda regionen för vargdomesticering.[5]

Med neolitiska revolutionen började människor bedriva selektiv avel, och skapade på så sätt hundraser. Nordamerikas indianer använde tidigt hunden som dragdjur.

Födoämnen, skötsel och vård

Trots att hunden ursprungligen var en typisk köttätare, har den som husdjur anpassats till att äta samma mat som människan och blivit en utpräglad allätare. Ständig tillgång till friskt dricksvatten är ett krav för hundens hälsa. Hundens lägerplats bör inte infekteras av parasiter. Ett tillfälligt bad är inte nödvändigt, men mycket nyttigt och hjälper till att hålla hunden i god kondition samt minskar den fräna lukt som kan orsakas av hundar som hålls inomhus. För unga hundar är en kraftig och närande diet av största vikt. Dels för att ge en kraftig kroppsbyggnad hos medelstora och stora hundraser och dels för att undvika valpsjukan. Teobromin som finns i kakaobönor och följaktligen i mörk choklad kan i större mängder orsaka livshotande teobrominförgiftning hos hundar. Det är inte nyttigt för en hund att äta födoämnen som innehåller mycket lök och salt heller.

I allmänhet är det viktigt för hundens psykiska utveckling att den får vistas så mycket som möjligt i människans sällskap. Det hjälper djuret även i intellektuellt avseende och skapar en bra relation mellan hunden och dess ägare.

Fortplantning och avel


Diande dalmatinervalpar.

Golden Retrievervalpar.
Tamhundens fortplantning är inte begränsad till någon viss årstid. Men de flesta tikar blir brunstiga (löper) två gånger om året, vanligen i januari eller februari och i juli eller augusti. När en tik och en hane parar sig med varandra, uppstår en förändring i hanens penis som gör att den sväller upp så att tiken och hanhunden inte kan skiljas från varandra, något som kallas för hängning. Parning kan ibland ske utan hängning, men då brukar tikens möjlighet att bli dräktig betraktas som mindre.

Efter dräktigheten, som tar omkring 63 dagar, föds valparna, som de första 9 till 12 dagarna är blinda. Antalet valpar är mycket växlande. Mindre hundraser får i allmänhet en till sju valpar medan medelstora eller stora raser föder mellan 6 och 10 valpar. I två fall (ett i Tyskland och ett i Danmark) var antalet valpar 26.[källa behövs] Eftersom tiken kan para sig flera gånger inför samma kull kan valparna i kullen härstamma från olika fäder. Detta syns tydligast när hanarna varit av olika ras.

Vid 6 veckors ålder kan valparna klara sig utan tikens mjölk. Bäst är att redan tidigare successivt vänja dem vid annan föda. Mjölktänderna börjar komma i 3:e eller 4:e veckan och ungefär vid 6 eller 7 veckors ålder är alla på plats. Tandömsningen sker i 3:e till 6:e månaden. Med fullbordad tandömsning upphör hundens valpperiod.

Mindre raser har vid denna tidpunkt nått sin slutliga storlek. Större raser växer ännu en tid, och de största blir fullstora först under tredje året. Könsmognaden inträder hos hanar vid en ålder av nio till elva månader. Tiken blir vanligtvis könsmogen under åttonde eller nionde månaden.

Små och medelstora hundar bör emellertid inte användas till avel innan de nått en ålder av 1½ eller 2 år och större raser inte förrän 3:e året, alltså tidigast vid den 3:e löpningen.[källa behövs] Under 3:e eller 4:e året når hunden sin högsta prestationsförmåga i detta avseende och redan under sjätte året förekommer ofta ett avtagande av rörlighet och krafter.[källa behövs] Hundens genomsnittsålder beräknas vanligen till 12 år, trots att några individer kan uppnå 18 års ålder och mer.[källa behövs] Den äldsta hunden blev 33 år gammal i Sverige.[källa behövs]

Hundens användningsområden


En svensk polishund.

En fårhund på jobbet.
Hundens användningsområden är många. Idag tränas det till och med upp hundar som kan upptäcka allvarliga sjukdomar, som cancer, på ett långt tidigare stadium än när något instrument kan klara den[källa behövs]. Man använder också så kallade epilepsihundar; hundar som är tränade att varna om ett kommande anfall, dämpa fallet om patienten faller, och till att hämta hjälp om det är nödvändigt[källa behövs].

Familjehundar

Familjehundar är hundar som är primärt rena familjehundar, som inte har någon annan uppgift än att glädja[6]. Studier har visat att hundens terapeutiska påverkan på människor ofta är positiv. Barn som växer upp med hund i huset lär sig ofta till exempel, att tidigare ta hänsyn.[6] Några hundar har också ibland övriga uppgifter som brukshundar, till exempel som jakthund eller slädhund.

Jakthundar

Jakthundar är hundar som används vid jakt. Det finns ett flertal olika hudraser som har avlats fram för olika former av jakt.

Brukshundar

En brukshund är en hund som per definition används för att lösa olika uppgifter. Den vanligaste brukshunden är en vakthund, hundar som aktivt eller passivt passar husdjur på bete eller bevakar egendom. Det finns både civila och offentliga tjänstehundar. En offentlig tjänstehund kan till exempel vara en militär tjänstehund eller en polishund tränade för olika uppgifter, exempelvis som patrullhund, narkotikahund eller en bombhund. En civil tjänstehund kan vara en servicehund med olika uppgifter, till exempel som ledarhund, hjälphund, vårdhund eller terapihund.

Hundsport

Hundsport är sportformer där hundar ingår som ett element. Lydnad, Spår, Sök, Skydd, Hundkapplöpning, agility,draghund, weight pulling

Utställning

Hundutställningar är populära bland personer som gillar att tävla om vem som har de mest rastypiska hundarna. En kvalificerad domare bedömer varje hund i hänvisning till en förhandsdefinierad och godkänd rasstandard för rasen, och därefter bedöms hundarna individuellt mot varandra könsvis, åldersvis, rasvis, gruppvis och till slut om vem som är den bästa utställningshunden på den aktuella utställningen.

Draghund


Hundkärra , 1904.
Draghundar används för transportändamål, vilket är fallet med slädhundar, men även andra typer av hundar har använts för sådant bruk. Sennenhundar användes för att dra kärror. Dalmatiner, liksom olika sorters gårdshundar nyttjades för att åtfölja ekipage med häst och vagn.

Draghundssport används som benämning för sådan hundsport vars ursprung kan hänföras till transportändamål. Weight pulling kan ses som en sådan hundsport.

Hundraser


Labrador retriever är en populär familjehund.
Begreppet hundras används för att beskriva så kallade rasrena hundar, det vill säga hundraser vars avelsarbete organiseras av en kennelklubb och där varje godkänd individ registreras och förses med en stamtavla som beskriver individens ursprung. Dock är nedanstående information av mer allmän karaktär och gäller oavsett ras eller blandningsförhållande.

Att välja en ras som passar

Att välja en ras som passar kan vara ett svårt val, om man först har bestämt sig för att bli hundägare. Dessvärre ser man allt för ofta att vissa familjer väljer fel ras, med resultatet att hunden antingen blir missanpassad i sin miljö, omplacerad eller i värsta fall avlivad. De allra flesta som skaffar sig hund ska primärt ha en familjehund, men det finns också de som letar efter den perfekta utställnings-, lydighets- eller brukshunden och som sätter sig extra bra in i blodslinjer, speciella kombinationer och avel. Några är också allergiska mot hundar, något som gör det svårt att ha hund.

Valets kval

När man väljer ras är det viktigt att välja en som passar till ens egen situation, miljö, aktivitets- och kompetensnivå. Det är således både dumt och naivt att tro att alla retriever är lydiga och välanpassade för att grannen har en sådan hund. Sådant kräver kunskap och träning. Likadeles är det dumt att välja en krävande och energisk vallhund om man ska ha en rolig, snäll och balanserad familjehund. Om man däremot är fårbonde och behöver en medhjälpare, är dessa raser ideala. Likadeles är det dumt att välja en typisk jakthund, som en fågelhund, om man inte själv är beredd att träna eller gå långa turer varje dag, även om man jagar ett par veckor på hösten. Energiska hundar passar bäst tillsammans med energiska människor, liksom bekväma hundar passar bäst med bekväma människor. Om man som bekväm människa önskar att skaffa hund för att få ett mer aktivt liv, bör man alltså först lägga om livsstilen och sedan skaffa sig en hund som passar efter att detta har lyckats. Mindre hundar brukar oftast behöva mindre motion, dock inte alla raser. Raser som framavlats som sällskapshundar är bättre anpassade till ett liv i lägenhet, med enstaka långpromenader. Det finns människor som vill ha lugn och ro omkring sig, då är det en misstag att välja en skällig hund. Hundraser som skäller mycket, som till exempel tax, chihuahua, foxterrier, cairnterrier, pekingese och i sådana fall måste vänjas av med att skälla för mycket redan från början, vilket kan vara en utmaning. Bäst att välja en tystylåten ras istället, som golden retriever, italiensk vinthund, vizsla, basenji, borzoi, japanese chin, chow chow, american water spaniel, clumber spaniel eller akita.[7][8]

Allergivänliga raser


Pudel räknas ofta som allergivänlig, men detta stöttas inte av forskningen.

Perro de agua español (Spansk vattenhund).
Hundallergi är egentligen bara ett annat ord för pälsdjursallergi. En sådan allergi kan utlösas av alla arter av pälsdjur, oavsett art, även alla typer hundar, eftersom alla pälsdjur producerar allergener - också nakenhundar och hundar med växande päls. Det finns således inga allergirena pälsdjur, men statistik visar på att färre reagerar på hundraser av typen ungersk puli, chinese crested dog /powder puff och pudel, men man vet inte varför, det kan vara en statistisk tillfällighet. Forskningen visar nämligen att det idag inte finns någon grund för att anta att det finns så kallade lågallergena hundraser eller pälsdjur. Det finns emellertid exempel på att några människor endast reagerar på bestämda pälsdjursarter eller raser, även om detta tillhör undantagen. Har man kraftig allergi kan man reagera på alla typer av pälsdjur, även i hus där det inte har bott sådana på flera månader.

Huvudallergenet, som heter Can d 1, har hittats i celler i hud, hår, serum, spott och urin hos alla pälsdjur. Det har också hittats hos alla undersökta hundraser, och det är lika stor variation på mängden allergen hos olika individer som det är mellan olika raser. Problemet är också i lika hög grad relaterat till andra arter, till exempel katter, marsvin, hästar, kor osv. Om djuren är små eller stora har heller ingen betydelse.

Om man fortfarande vill skaffa sig en hund, eller ett annat pälsdjur, bör man välja ett djur som har tät växande päls och därför måste trimmas eller klippas regelbundet. Ett sådant djur är att föredra framför ett djur som har vinterpäls eller helt saknar hår, men bara om de kan badas ofta. Exempel på sådana pälsdjur är hundraser som portugisisk vattenhund, bichon frisé, old english sheepdog, pudel, irish softcoated wheaten terrier, tibetansk terrier, chinese crested dog, powder puff och ungersk puli och komondor med flera. Det är emellertid en förutsättning att djuret badas ofta, kanske flera gånger i veckan, för också sådana djur har allergener som kan (kommer att) utlösa allergiska reaktioner.

Vilka hundraser man "tål" varierar också beroende på hur allergisk just Du är. Många tycker att det är en bra idé att åka hem till uppfödare av de raser som är allergivänliga, dock kan man reagera ändå; uppfödaren kan ha andra raser, eller många hundar, och då kan man få en allergisk reaktion.

Svenska hundraser


Jämthund godkändes som egen ras 1946, dessförinnan sågs den som en otypiskt stor gråhund.[9]
Det finns elva svenska hundraser[9] som är erkända av SKK. Tio av dessa är erkända i alla nordiska länder och åtta är internationellt erkända av den internationella kennelfederationen Fédération Cynologique Internationale (FCI). För en tolfte ras, dansk/svensk gårdshund, delas ansvaret mellan Sverige och Danmark, denna ras är interimerkänd av FCI sedan 2008. Härutöver har Nordisk Kennelunion (NKU) gemensamt avelsansvar för samojedhunden med ursprung i norra Ryssland och Sibirien. Även gråhund har räknats som svensk men 1981 slogs denna ihop med norsk älghund, grå. Tidigare har den danska strellufstövaren slagits samman med den svenska drevern. Dessutom bedrivs avel med hedehund, en nordlig jaktspets (älghund) som inte är en erkänd ras. En utdöd svensk hundras är dalbohunden som var av molossertyp. Som Sveriges nationalras räknas hamiltonstövaren som är namngiven efter SKK:s förste ordförande Adolf Patrik Hamilton[9].


Hamiltonstövare , Sveriges nationalras.
Dansk/svensk gårdshund (gårdshund / pinscher, FCI)
Drever (drivande hund, FCI)
Gotlandsstövare (drivande hund / stövare, endast SKK)
Hamiltonstövare (drivande hund / stövare, FCI)
Hälleforshund (älghund / nordlig jaktspets, NKU)
Jämthund (älghund / nordlig jaktspets, FCI)
Norrbottenspets (skällande fågelhund / nordlig jaktspets, FCI)
Schillerstövare (drivande hund / stövare, FCI)
Smålandsstövare (drivande hund / stövare, FCI)
Svensk lapphund (vallande spets, FCI)
Svensk vit älghund (älghund / nordlig jaktspets, NKU)
Västgötaspets (gårdshund / vallande spets, FCI)
Förbjudna hundraser


Pitbullterrier klassas normalt som en kamphundsras.
I många länder har flera hundraser på senare år blivit förbjudna att hålla, eftersom lokala myndigheter räknar hundarna som speciellt farliga. Förbudet omfattar många så kallade kamphundar, men många länder har också förbjudit blandningshundar där förbjudna raser eller varg ingår.[källa behövs]

Grundanledningen till förbudet var att det började växa fram olagliga etableringar av kamphundsmiljöer, där reguljära hundkamper arrangerades för pengarnas (vadslagning) eller för nöjes skull. Dessa miljöer etablerades först i USA, men spred sig sedan snabbt till andra länder i den industrialiserade världen.

Övrigt och kuriosa

Kanarieöarna har fått sitt namn efter det latinska ordet canis, och betyder alltså hundöarna. "Hundarna" det syftas på tros dock vara sälar ("sjöhundar").[källa behövs]
Den snabbaste hundrasen, greyhound, kan på kortare sträckor springa 70 kilometer i timmen.[10]
Galleri


Engelsk bulldogg

 

Alaskan malamute

 

Beagle

 

Chihuahua

 

Chow chow

 

Dalmatiner

 

Schäfer

 

Golden retriever

 

Pudel

 

Dvärgschnauzer

 

Dvärgpinscher

 

Västgötaspets

 

Puli

 

Tibetansk terrier

 

Kinesisk nakenhund

Se även

Hundens historia
Hundsjukdomar
Gruppindelning av hundraser
Lista över berömda hundar
Källor

Artikeln är delvis en översättning från Wikipedia på norska (bokmål)
Hunden i Nordisk familjebok (andra upplagan, 1909)
Noter

